//CounterInput: 4-bit input to determine what mode to run
//CounterEnable: 1-bit input to determine if counter is on (Only on if coin is inserted)


module Counter_Main(CounterInput, CounterEnable, Clk, nReset, S0, S1, S2);
